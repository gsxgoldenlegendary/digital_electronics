`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 26.11.2021 17:59:13
// Design Name:
// Module Name: VRAM
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module VRAM(input [14:0]raddr,
            input [14:0]waddr,
            [11:0]wdata,
            we,
            output [11:0]rdata);
            
endmodule
